.title KiCad schematic
.model __Q1 NPN
.model __Q2 NPN
.model __Q4 NPN
.model __Q3 NPN
.model __Q7 NPN
.model __Q6 NPN
.model __Q5 PNP
R37 GND /SPI_MUX_SEL 10k
U7 __U7
C17 +3.3V GND 1u
C8 Net-_U8-XTAL2_ GND 15p
Y1 __Y1
C13 Net-_U8-XTAL1_ GND 15p
C10 Net-_U8-AREF_ GND 10u
C14 Net-_U8-AREF_ GND 100n
SW3 __SW3
J3 __J3
C12 +3.3V GND 100n
C9 +3.3V GND 100n
FID2 __FID2
FID3 __FID3
FID4 __FID4
H4 __H4
FID1 __FID1
H1 __H1
H3 __H3
H2 __H2
R5 Net-_J2-DAT1_ /CDAT1 100
R6 Net-_J2-DAT0_ /CDAT0 100
R7 /CCLK Net-_J2-CLK_ 100
R9 /CDAT3 Net-_J2-CD/DAT3_ 100
R8 /CCMD Net-_J2-CMD_ 100
R10 /CDAT2 Net-_J2-DAT2_ 100
J2 __J2
C3 /VTM GND 100n
R17 /LED_U3 Net-_Q2-B_ 1k
R25 Net-_D4-K_ Net-_Q2-C_ 270
R12 Net-_U1-KVBUS_ GND 1k
R11 VBUS Net-_U1-KVBUS_ 1k
C1 +3.3V GND 100n
C2 /CLDO GND 100n
R1 /RREF GND 6.19k
R2 GND /mode 10k
U1 __U1
JP1 __JP1
R15 +3.3V Net-_U3-DCNF0_ 1k
R18 Net-_D2-K_ /UART_RX_LED 270
D1 __D1
R14 Net-_D1-K_ /UART_TX_LED 270
C7 +3.3V GND 100n
U4 __U4
R35 SCL_I2C +3.3V 1k
TP2 __TP2
R27 Net-_U4-_RESET_ +3.3V 1k
R34 SDA_I2C +3.3V 1k
R20 /SDA_MCU +3.3V 1k
R19 /SCL_MCU +3.3V 1k
R21 /SCL_USB +3.3V 1k
R23 /SDA_USB +3.3V 1k
JP2 __JP2
R32 Net-_U3-DM_ USB_FTDI_D- 33
U3 __U3
TP1 __TP1
R26 VBUS Net-_U3-VBUS_DET_ 5.1k
R13 +3.3V Net-_U3-DCNF1_ 1k
D2 __D2
C5 +3.3V GND 100n
R31 Net-_U3-DP_ USB_FTDI_D+ 33
C6 +3.3V GND 4.7u
R36 RST# Net-_JP2-A_ 100
R39 /EXT_I2C_EN +3.3V 10k
U10 __U10
J4 __J4
U11 __U11
Y2 __Y2
C18 +3.3V GND 100n
C19 Net-_U11-VBAT_ GND 100n
U8 __U8
C11 /RST#_P RST# 4.7u
R38 /RST#_P +3.3V 10k
C15 +3.3V GND 100n
C16 +3.3V GND 100n
U5 __U5
U6 __U6
U9 __U9
J1 __J1
R24 Net-_D3-K_ Net-_Q1-C_ 270
R22 +3.3V /BTN_USER_A 10k
SW1 __SW1
D3 __D3
R16 /LED_U1 Net-_Q1-B_ 1k
Q1 Net-_Q1-B_ GND Net-_Q1-C_ __Q1
Q2 Net-_Q2-B_ GND Net-_Q2-C_ __Q2
D4 __D4
R29 /buzzer Net-_Q4-B_ 1k
Q4 Net-_Q4-B_ GND Net-_BZ1-+_ __Q4
Q3 Net-_Q3-B_ GND Net-_Q3-C_ __Q3
R30 +3.3V /BTN_USER_B 10k
SW2 __SW2
BZ1 __BZ1
R33 Net-_D5-K_ Net-_Q3-C_ 270
D5 __D5
R28 /LED_U2 Net-_Q3-B_ 1k
R4 GND Net-_J1-CC1_ 5.1k
R3 GND Net-_J1-CC2_ 5.1k
U2 __U2
C4 VBUS GND 1n
NT1 __NT1
R52 Net-_BT1A--_ GND 0R01 75PPM
NT2 __NT2
D11 __D11
D12 __D12
D10 __D10
D8 __D8
D9 __D9
D15 __D15
D14 __D14
D13 __D13
R60 Net-_D15-K_ /liion/H 270
R53 Net-_D8-K_ /liion/A 270
C33 +3.3V GND 100n
U14 __U14
R54 Net-_D9-K_ /liion/B 270
R55 Net-_D10-K_ /liion/C 270
R57 Net-_D12-K_ /liion/E 270
R56 Net-_D11-K_ /liion/D 270
R59 Net-_D14-K_ /liion/G 270
R58 Net-_D13-K_ /liion/F 270
F5 __F5
F4 __F4
BT1 __BT1
F2 __F2
F3 __F3
BT2 __BT2
F1 __F1
C21 Net-_U13-PMID_ GND 100n
C20 Net-_U13-PMID_ GND 10u
R50 Net-_U13-TS_BIAS_ Net-_U13-TS_ 5.3k
R47 Net-_U13-ILIM_ GND 2.49k
C24 Net-_U13-ILIM_ GND 1u
C30 +BATT GND 10u
TH2 __TH2
C32 Net-_U13-REGN_ GND 4.7u
R51 Net-_U13-TS_ Net-_R51-Pad2_ 31.1k
U13 __U13
L1 Net-_U13-SW_ +VSW 1uH - DFE252012P-1R0M=P2
C29 Net-_U13-SW_ Net-_U13-BTST_ 47n
C31 +VSW GND 22u
R49 /liion/GAUGE_SRN Net-_U12-SRN_ 100
C26 Net-_U12-SRP_ GND 100n
C27 Net-_U12-SRN_ GND 100n
C23 Net-_U12-SRP_ Net-_U12-SRN_ 100n
Q7 Net-_Q7-B_ GND Net-_Q7-C_ __Q7
R42 /liion/CH_PG Net-_Q7-B_ 1k
R41 /liion/CH_STAT Net-_Q6-B_ 1k
Q6 Net-_Q6-B_ GND Net-_Q6-C_ __Q6
D6 __D6
R45 Net-_D6-K_ Net-_Q6-C_ 270
D7 __D7
R46 Net-_D7-K_ Net-_Q7-C_ 270
SW4 __SW4
C28 Net-_U12-REG25_ GND 1u
C25 /liion/Battery+ GND 3.3n
TH1 __TH1
R48 /liion/GAUGE_SRP Net-_U12-SRP_ 100
C22 +3.3V GND 100n
U12 __U12
R44 GND /liion/GAUGE_BTN_IN 1k
R40 /liion/CH_BTN Net-_Q5-B_ 510
Q5 Net-_Q5-B_ +3.3V Net-_Q5-C_ __Q5
R43 /liion/GAUGE_BTN_IN Net-_Q5-C_ 270
U15 __U15
L2 Net-_U15-LX1_ Net-_U15-LX2_ 1uH - DFE252012P-1R0M=P2
C34 +VSW GND 22u
R62 GND EXT_PWR_5v_EN 1k
C36 +VSW GND 22u
R63 /sw_source/5v_mod +VSW 1k
JP6 __JP6
L4 Net-_U17-LX1_ Net-_U17-LX2_ 1uH - DFE252012P-1R0M=P2
C39 5v_EXT GND 47u
R70 5v_EXT /sw_source/5v_FB 806k
R71 /sw_source/5v_FB GND 91k
U17 __U17
C42 5v_EXT GND 10u
C46 3v3_SD GND 100n
C45 3v3_SD GND 10u
C44 Net-_U18-CT_ GND 1n
L5 Net-_L5-Pad1_ 3v3_SD 100u
U18 __U18
C43 +3.3V GND 1u
C41 3v3_EXT GND 10u
C38 3v3_EXT GND 47u
R68 3v3_EXT /sw_source/3v3_FB 511k
R69 /sw_source/3v3_FB GND 91k
U16 __U16
L3 Net-_U16-LX1_ Net-_U16-LX2_ 1uH - DFE252012P-1R0M=P2
C35 +VSW GND 22u
R64 /sw_source/3v3_mod +VSW 1k
R61 GND EXT_PWR_3v3_EN 1k
JP5 __JP5
JP7 __JP7
R65 /sw_source/3v3i_mod +VSW 1k
JP4 __JP4
JP3 __JP3
R66 +3.3V /sw_source/3v3i_FB 511k
C37 +3.3V GND 47u
R67 /sw_source/3v3i_FB GND 91k
C40 +3.3V GND 10u
.end
